** Profile: "SCHEMATIC1-simulare_frecv"  [ C:\Users\TEO\Desktop\P1_2024_431A_CatrinescuTeodora_PAI_nr24_Orcad\pai\pai-pspicefiles\schematic1\simulare_frecv.sim ] 

** Creating circuit file "simulare_frecv.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 10 1 10000k
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
